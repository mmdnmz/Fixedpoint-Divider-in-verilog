module sub (input [10:0] a, b, output [10:0] c);

  assign c = a - b;
endmodule
